(* Require Import OrderedType Relations. *)
(* Require FSets.OrderedType FSets.OrderedTypeAlt. *)

(* (** This file contains conversion facilities between typeclass-based *)
(*    ordered types and module-bases ordered types. *) *)

(* (** * From typeclasses to modules *) *)

(* (** ** Constructing an [OrderedType] module *)

(*    This functor creates an [FSets.OrderedType.OrderedType] module for a  *)
(*    type [t] given an [OrderedType t] instance. The input signature [S] of  *)
(*    the functor is just a module packing a type and an instance together. *)

(*    Note that using this functor is one way of ensuring by construction that *)
(*    the computational and specification parts of the [compare] function in *)
(*    the [OrderedType] module are adequately separated. *)
(*    *) *)
(* Module Type S. *)
(*   Parameter t : Type. *)
(*   Instance Ht : OrderedType t. *)
(* End S. *)

(* Module OT_to_FOT (Import X : S) <: OrderedType.OrderedType. *)
(*   Definition t := t. *)

(*   Definition eq : relation t := _eq. *)
(*   Definition lt : relation t := _lt. *)

(*   Definition eq_refl : forall (x : t), eq x x := reflexivity. *)
(*   Definition eq_sym : forall (x y : t), eq x y -> eq y x := symmetry. *)
(*   Definition eq_trans : forall (x y z : t), eq x y -> eq y z -> eq x z :=  *)
(*     transitivity. *)

(*   Definition lt_not_eq : forall (x y : t), lt x y -> ~eq x y := lt_not_eq. *)
(*   Definition lt_trans : forall (x y z : t), lt x y -> lt y z -> lt x z :=  *)
(*     transitivity. *)

(*   Definition compare_1 : forall x y, x =?= y = Eq -> eq x y. *)
(*   Proof. intros x y; destruct (compare_dec x y); intuition discriminate. Qed. *)
(*   Definition compare_2 : forall x y, x =?= y = Lt -> lt x y. *)
(*   Proof. intros x y; destruct (compare_dec x y); intuition discriminate. Qed. *)
(*   Definition compare_3 : forall x y, x =?= y = Gt -> lt y x. *)
(*   Proof. intros x y; destruct (compare_dec x y); intuition discriminate. Qed. *)
(*   Definition compare : forall x y, OrderedType.Compare lt eq x y. *)
(*   Proof. *)
(*     intros x y; case_eq (x =?= y); intro Hcomp. *)
(*     constructor 2; exact (compare_1 _ _ Hcomp). *)
(*     constructor 1; exact (compare_2 _ _ Hcomp). *)
(*     constructor 3. exact (compare_3 _ _ Hcomp). *)
(*   Defined. *)

(*   Definition eq_dec : forall x y, {eq x y} + {~(eq x y)}. *)
(*   Proof. *)
(*     intros; case_eq (x =?= y); intro Hcomp. *)
(*     left; exact (compare_1 _ _ Hcomp). *)
(*     right; apply lt_not_eq; exact (compare_2 _ _ Hcomp). *)
(*     right; apply gt_not_eq; exact (compare_3 _ _ Hcomp). *)
(*   Defined. *)
(* End OT_to_FOT. *)

(* (** ** Constructing an [OrderedTypeAlt] module *)

(*    This functor creates an [FSets.OrderedType.OrderedTypeAlt] module  *)
(*    for a type [t] given an [OrderedType t] instance.  *)

(*    Make sure you use this functor instead of combining the functor [OT_to_FOT] *)
(*    above and the functor [OrderedType_to_Alt] from the standard library to  *)
(*    avoid loss of performance in the comparison function. *)
(*    *) *)
(* Module OT_to_FOT_Alt (Import X : S) <: OrderedTypeAlt.OrderedTypeAlt. *)
(*   Definition t := t. *)

(*   Definition compare (x y : t) := x =?= y. *)

(*   Property compare_sym : forall x y, (compare y x) = CompOpp (compare x y). *)
(*   Proof. *)
(*     intros; unfold compare; destruct (compare_dec x y);  *)
(*       destruct (compare_dec y x); order. *)
(*   Qed. *)

(*   Property compare_trans : *)
(*     forall c x y z, compare x y = c -> compare y z = c -> compare x z = c. *)
(*   Proof. *)
(*     intros; unfold compare in *;  *)
(*       destruct (compare_dec x y); destruct (compare_dec y z); *)
(*         destruct (compare_dec x z); auto; order; congruence. *)
(*   Qed. *)
(* End OT_to_FOT_Alt. *)

(* (** * From modules to typeclasses *) *)

(* (** ** Constructing an instance from an [OrderedType] module *)

(*    This functor creates an [OrderedType] instance given a *)
(*    [FSets.OrderedType.OrderedType] module. *)

(*    Use with caution because, depending on the design of the original *)
(*    [compare] function, the comparison function in the resulting instance *)
(*    may compute 'proofs' that are discarded in the end.     *)
(*    *) *)
(* Module FOT_to_OT (Import X : OrderedType.OrderedType). *)
(*   Section ForInstances. *)
(*     Instance eq_Equivalence : Equivalence eq := { *)
(*       Equivalence_Reflexive := eq_refl; *)
(*       Equivalence_Symmetric := eq_sym; *)
(*       Equivalence_Transitive := eq_trans *)
(*     }. *)

(*     Instance lt_StrictOrder : StrictOrder lt eq := { *)
(*       StrictOrder_Irreflexive := lt_not_eq; *)
(*       StrictOrder_Transitive := lt_trans *)
(*     }. *)
(*   End ForInstances. *)

(*   Definition cmp (x y : X.t) := *)
(*     match compare x y with *)
(*       | OrderedType.LT _ => Lt *)
(*       | OrderedType.EQ _ => Eq *)
(*       | OrderedType.GT _ => Gt *)
(*     end. *)
(*   Program Instance t_OT : OrderedType X.t := { *)
(*     _eq := eq; *)
(*     _lt := lt; *)
(*     OT_Equivalence := eq_Equivalence; *)
(*     OT_StrictOrder := lt_StrictOrder; *)
(*     _cmp := cmp *)
(*   }. *)
(*   Next Obligation. *)
(*     unfold cmp; destruct (compare x y); constructor; auto. *)
(*   Qed. *)
(* End FOT_to_OT. *)

(* (** ** Constructing an instance from an [OrderedTypeAlt] module  *)

(*    This functor creates an [OrderedType] instance given a *)
(*    [FSets.OrderedType.OrderedTypeAlt] module. *)
(*    *) *)
(* Module FOT_Alt_to_OT (Import X : OrderedTypeAlt.OrderedTypeAlt). *)
(*   Definition eq (x y : t) := x ?= y = Eq. *)
(*   Definition lt (x y : t) := x ?= y = Lt. *)

(*   Section ForInstances. *)
(*     Program Instance eq_Equivalence : Equivalence eq. *)
(*     Next Obligation. (* reflexivity *) *)
(*       intro x; unfold eq. *)
(*       assert (H := compare_sym x x); destruct (x ?= x); auto; discriminate. *)
(*     Qed. *)
(*     Next Obligation. (* symmetry *) *)
(*       intros x y; unfold eq. *)
(*       generalize (compare_sym x y); assert (H := fun c => compare_trans c x y x); *)
(*         destruct (x ?= y); destruct (y ?= x); auto; simpl; intros; discriminate. *)
(*     Qed. *)
(*     Next Obligation. (* transitivity *) *)
(*       intros x y z; unfold eq. *)
(*       exact (compare_trans Eq x y z). *)
(*     Qed. *)

(*     Program Instance lt_StrictOrder : StrictOrder lt eq := { *)
(*       StrictOrder_Irreflexive := _; *)
(*       StrictOrder_Transitive := _ *)
(*     }. *)
(*     Next Obligation. (* transitivity *) *)
(*       intros x y z; unfold lt. *)
(*       exact (compare_trans Lt x y z). *)
(*     Qed. *)
(*     Next Obligation. (* irreflexivity *) *)
(*       intros abs; compute in abs; unfold lt in H; destruct (x ?= y); congruence. *)
(*     Qed. *)
(*   End ForInstances. *)

(*   Definition cmp (x y : X.t) := x ?= y. *)
(*   Program Instance t_OT : OrderedType X.t := { *)
(*     _eq := eq; *)
(*     _lt := lt; *)
(*     OT_Equivalence := eq_Equivalence; *)
(*     OT_StrictOrder := lt_StrictOrder; *)
(*     _cmp := cmp *)
(*   }. *)
(*   Next Obligation. *)
(*     unfold cmp; case_eq (x ?= y); constructor; auto. *)
(*     unfold lt; rewrite (compare_sym x y); rewrite H; auto. *)
(*   Qed. *)
(* End FOT_Alt_to_OT. *)
